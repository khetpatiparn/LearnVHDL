library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity T14_CaseWhenTb is
end entity;
	
architecture sim of T14_CaseWhenTb is
	
begin
	process is
	begin
	
	end process;
	

end architecture;