library ieee;
use ieee.std_logic_1164.all;

entity T17_ClockProcessTb is
end entity;

architecture sim of T17_ClockProcessTbr is

	
begin

	process is
	begin

	end process;

end architecture;